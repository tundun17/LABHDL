module Dem (
    input 
);
    
endmodule